

package my_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh";
    `include "adder_transaction.sv";
    `include "uvm_driver.sv";
    `include "uvm_sequencer.sv";
    `include "uvm_agent.sv";
    `include "uvm_sequence.sv";
    `include "uvm_sequence2.sv";
    `include "seq_of_sequences.sv";
    `include "uvm_envt.sv";
    `include "uvm_test.sv";
    
    

endpackage